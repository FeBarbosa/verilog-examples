module test_adder(a, b, s, cin, cout);
	input a;
	input b;
	input cin;
	
	output s;
	output cout;

	assign s =  a ^ b ^ cin;
	assign cout =  a & b | a & cin | b & cin;
endmodule // test_adder
